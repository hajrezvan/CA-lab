--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   22:12:32 03/07/2022
-- Design Name:   
-- Module Name:   D:/ISE/experiment_1/experiment_3/up_tb.vhd
-- Project Name:  experiment_3
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: up
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY up_tb IS
END up_tb;
 
ARCHITECTURE behavior OF up_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT up
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         q : INOUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';

	--BiDirs
   signal q : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: up PORT MAP (
          clk => clk,
          reset => reset,
          q => q
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		reset <= '1';
      -- hold reset state for 100 ns.
      wait for 50 ns;
		reset <= '0';
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
		wait for 50 ns;
      wait for 50 ns;

      wait;
   end process;

END;
